`timescale 1ns / 1ps

module program_memory (
    input clk,
    input [31:0] byte_address,
    input write_enable,         
    input [31:0] write_data, 
    output logic [31:0] read_data
    // output logic [31:0] curr_read_data,
    // output logic [31:0] next_read_data
);

    logic [31:0] ram [0:255];
    logic [7:0] word_address;
    
    
    assign word_address = byte_address[9:2];
    
    
    // initial begin
        // $readmemb("instruction_mem.mem", ram);  the reading process is not functional
        // test for LW,ADD instructions, temporarily
        // ram[0] = 32'b00000000001100000000000110000011; // LW x1, 3(x0)
        // ram[1] = 32'b00000000011000000000001010000011; // LW x2, 6(x0)
        // ram[2] = 32'b00000000000000000000000000010011; // NOP
        // ram[3] = 32'b00000000001000001000000110110011; // ADD x3,x1,x2
        // ram[4] = 32'b00000000000000000000000000010011; // NOP
        // ram[5] = 32'b00000000001100000010001000100011; // SW x3,8(x0)

        // test for ADDI, ADD instructions 
        // funct 7 rs2 rs1 funct3 rd opcode , solved related bugs.
        //ram[0] = 32'b00000000_00000_00000_000_00000_0010011; //nop
        //ram[1] = 32'b00000000_00001_00000_000_00001_0010011; // (ADDI x1, x0, 1)
        //ram[2] = 32'b00000000_00010_00000_000_00010_0010011; //(ADDI x2, x0, 2)
        //ram[3] = 32'b00000000_00011_00000_000_00011_0010011; // (ADDI x3, x0, 3)
        //ram[4] = 32'b00000000_00100_00001_000_00100_0010011; // (ADDI x4, x1, 4)
        //ram[5] = 32'b00000000_00010_00011_000_00101_0110011; //(ADD X5,X1,X2)
        //ram[6] = 32'b00000000_00000000_00010001_00010001; // end transition

        // test for branch with initial taken and not taken, test flush, jal, jalr
        // ram[0] = 32'b0000000_00011_00000_000_00010_0010011; // ADDI x2, x0, 3
        // ram[1] = 32'b0000000_00101_00000_000_00001_0010011; //ADDI x1, x0, 5      
        // // imm[12] = 0; +imm[10:5] = 000000; +rs2 +rs1 +funt3 +im[4:1] = 1010 + imm[11] = 0 + opcode
        // // 20 = 0_0000_0001_0100
        // ram[2] = 32'b0000000_00001_00010_000_1010_0_1100011;// beq x2,x1 offset is 20
        // ram[3] = 32'b0000000_00001_00000_000_00100_0010011; // (addi x4,x0,1)
        // ram[4] = 32'b0000000_00001_00010_000_00010_0010011; // (addi x2, x2, 1 predition fail) 
        // ram[5] = 32'b0000000_00000_00000_000_00000_0010011; // nop     
        // ram[6] = 32'b1_1111111000_1_11111111_00000_1101111; // jal pc-16
        // // im[20]=1,im[10:1]=11111111000,im[11]=1,im[19:12]=11111111;rd=00000,opcode=1101111;
        // // -16 = 13'b111111111111111110000
        // ram[7] = 32'b0000000_01111_00000_000_00011_0010011; //label: addi x3, x0, 15)
        // ram[8] = 32'b0000000_00110_00000_000_01000_0010011; //x8 =6;
        // ram[8] = 32'b0000000_00000_00000_000_00000_0010011; // (end: nop)*/


        // ram[0] = 32'h0020_0093; // addi x1, x0, 2
        // ram[1] = 32'h0593_4529; // c.li x10, 10; then half of addi x11, x0, 5
        // ram[2] = 32'h061d_0050; // half of addi x11, x0, 5; then c.addi x12, 7
        // ram[3] = 32'h0030_0693; // addi x13, x0, 3
        // ram[4] = 32'h458d_9506; // c.add x10, x1; then c.li x11, 3
        // ram[5] = 32'h862a_8d0d; // c.sub x10, x11; then c.mv x12, x10
        // ram[6] = 32'h8909_8e69; // c.and x12, x10; then c.andi x10, 2
        // ram[7] = 32'h8d35_8e49; // c.or x12, x10; then c.xor x10, x13
        // ram[8] = 32'h0592_6595; // c.lui x11, 5; then c.slli x11, 4
        // ram[9] = 32'h0713_8591; // c.srai x11, 4; then half of addi x14, x0, -1
        // ram[10] = 32'h8311_fff0; // half of addi x14, x0, -1; then c.srli x14, 4
        // ram[11] = 32'h42d0_c2cc; // c.sw x11, 4(x13), then c.lw x12, 4(x13)

        // test 3
        // ram[0] = 32'b11111110110111001100101000110111;
        // ram[1] = 32'b00000000000010100000101000010011;
        // ram[2] = 32'b10101001100010100000101000010011;
        // ram[3] = 32'b00000000011010101000101010010011;
        // ram[4] = 32'b00000001010010101000101100110011;
        // ram[5] = 32'b01000001011010100000101110110011;
        // ram[6] = 32'b00000000000010111000110000110011;
        // ram[7] = 32'b01000001100000000000110000110011;
        // ram[8] = 32'b00000000000000000000000000010011;
        // ram[9] = 32'b00000000000000000000000000010011;

        // // test 4
        // ram[0] = 32'b00000000000100000000010100010011;
        // ram[1] = 32'b00000000100000000000000011101111;
        // ram[2] = 32'b00000101010000000000000011101111;
        // ram[3] = 32'b00000000000111110010000000100011;
        // ram[4] = 32'b00000000101011110010001000100011;
        // ram[5] = 32'b00000000100011110000111100010011;
        // ram[6] = 32'b11111111111101010000010110010011;
        // ram[7] = 32'b00000000000000000000000000010011;
        // ram[8] = 32'b00000000000000000000000000010011;
        // ram[9] = 32'b00000000000001011101100001100011;
        // ram[10] = 32'b00000000000000000000010100010011;
        // ram[11] = 32'b11111111100011110000111100010011;
        // ram[12] = 32'b00000000000000001000000001100111;
        // ram[13] = 32'b11111111111101010000010100010011;
        // ram[14] = 32'b11111101010111111111000011101111;
        // ram[15] = 32'b00000000000001010000101000010011;
        // ram[16] = 32'b11111111100011110000111100010011;
        // ram[17] = 32'b00000000010011110010010100000011;
        // ram[18] = 32'b00000000000011110010000010000011;
        // ram[19] = 32'b00000001010001010000010100110011;
        // ram[20] = 32'b00000000000000000000000000010011;
        // ram[21] = 32'b00000000000000000000000000010011;
        // ram[22] = 32'b00000000000000001000000001100111;
        // ram[23] = 32'b00000000000000000000000000010011;
        // ram[24] = 32'b00000000000000000000000000010011;

        // // test 5
        // ram[0] = 32'b10101001100001110110000010110111;
        // ram[1] = 32'b01010100001100001000000010010011;
        // ram[2] = 32'b00000000000100000010000000100011;
        // ram[3] = 32'b00000000000000000000000100000011;
        // ram[4] = 32'b00000000000100000000000110000011;
        // ram[5] = 32'b00000000001000000000001000000011;
        // ram[6] = 32'b00000000001100000000001010000011;
        // ram[7] = 32'b00000000000000000001001110000011;
        // ram[8] = 32'b00000000001000000001010000000011;
        // ram[9] = 32'b00000000000000000010010100000011;
        // ram[10] = 32'b00000000010000000010010110000011;
        // ram[11] = 32'b00000000000000000000000000010011;
        // ram[12] = 32'b00000000000000000000000000010011;
        // ram[13] = 32'b00000000000000000000000000010011;


        // // test 6
        // ram[0] = 32'h0000_0613;  // addi x12, x0, 0
        // ram[1] = 32'h0030_0693;  // addi x13, x0, 3
        // ram[2] = 32'h0000_0713;  // addi x14, x0, 0
        // ram[3] = 32'h0813_4785;  // c.li x15, 1; then half of addi x16, x0, 1
        // ram[4] = 32'h0001_0010;  // half of addi x16, x0, 1; then c.nop
        // // store_loop
        // ram[5] = 32'h0016_0613;  // addi x12, x12, 1
        // ram[6] = 32'h00f7_2023;  // sw x15, 0(x14)
        // ram[7] = 32'h0107_97b3;  // sll x15, x15, x16
        // ram[8] = 32'h0047_0713;  // addi x14, x14, 4
        // ram[9] = 32'hfed6_48e3;  // blt x12, x13, store_loop

        // ram[10] = 32'h0000_0613;  // addi x12, x0, 0
        // ram[11] = 32'h0000_0713;  // addi x14, x0, 0
        // ram[12] = 32'h0000_0413;  // addi x8, x0, 0
        // ram[13] = 32'hfff6_8693;  // addi x13, x13, -1
        // // load_loop
        // ram[14] = 32'h2783_0605;  // c.addi x12, 1; then half of lw x15, 0(x14)
        // ram[15] = 32'h0713_0007;  // half of lw x15, 0(x14); then addi x14, x14, 4
        // ram[16] = 32'h8c3d_0047;  // half of addi x14, x14, 4; then c.xor x8, x15
        // ram[17] = 32'hfec6_dae3;  // bge x13, x12, load_loop
        // ram[18] = 32'h0000_0013;  // nop

        // test 7
        // ram[0] = 32'h0000_0093; // addi x1, x0, 0
        // ram[1] = 32'h448d_4415; // c.li x8, 5; then c.li x9 3
        // ram[2] = 32'h14f9_94a2; // c.add x9, x8; then c.addi x9, -2
        // ram[3] = 32'h8c89_453d; // c.li x10, 15; then c.sub x9, x10
        // ram[4] = 32'h8085_0506; // c.slli x10, 1; then c.srli x9, 1
        // ram[5] = 32'hc388_4781; // c.li x15, 0; then c.sw x10, 0(x15)
        // ram[6] = 32'h0791_c3c4; // c.sw x9, 4(x15); then c.addi x15, 4
        // ram[7] = 32'ha603_438c; // c.lw x11, 0(x15); then low half of lw x12, -4(x15)
        // ram[8] = 32'h86aa_ffc7; // high half of lw x12, -4(x15); then c.mv x13, x10
        // ram[9] = 32'hc699_8e91; // c.sub x13, x12; then c.beqz x13, l
        // ram[10] = 32'h0010_8093; // addi x1, x1, 1
        // ram[11] = 32'h0010_8093; // addi x1, x1, 1
        // ram[12] = 32'h0010_8093; // addi x1, x1, 1
        // ram[13] = 32'h1230_8093; // l: addi x1, x1, 0x123
        // ram[14] = 32'h0000_0013; // nop
        // ram[15] = 32'h0000_0013; // nop

        // // test 8
        // ram[0] = 32'h8000_0437; // lui x8, 0x8000
        // ram[1] = 32'h0004_0413; // addi x8, x8, 0
        // ram[2] = 32'hffff_f4b7; // lui x9, 0xffff
        // ram[3] = 32'h0001_44bd; // c.li x9, 15; then c.nop
        // // loop:
        // ram[4] = 32'hfff4_8493; // addi x9, x9, -1
        // ram[5] = 32'h0013_8405; // c.srai x8, 1; then low half of nop
        // ram[6] = 32'hf8fd_0000; // high half of nop; then c.bnez x9, loop
        // ram[7] = 32'h0000_0013; // nop
        // ram[8] = 32'h0000_0013; // nop

        // // benchmark
        // ram[0]  = 32'h00a0_0513; // 0000_0000_1010_0000_0000_0101_0001_0011
        // ram[1]  = 32'h00c0_00ef; // 0000_0000_1100_0000_0000_0000_1110_1111
        // ram[2]  = 32'h0000_0013; // 0000_0000_0000_0000_0000_0000_0001_0011
        // ram[3]  = 32'h08c0_006f; // 0000_0111_1100_0000_0000_0110_0110_1111
        // // MATRIX_SUM_OF_PRODUCTS
        // ram[4]  = 32'h0000_0693; // 0000_0000_0000_0000_0000_0110_1001_0011
        // ram[5]  = 32'h0000_0313; // 0000_0000_0000_0000_0000_0011_0001_0011
        // ram[6]  = 32'h0000_0213; // 0000_0000_0000_0000_0000_0100_0001_0011
        // ram[7]  = 32'h0000_0013; // 0000_0000_0000_0000_0000_0000_0001_0011
        // // LOOP_I
        // ram[8]  = 32'h06a1_8a63; // 0000_0110_1010_0011_0000_0100_0110_0011
        // ram[9]  = 32'h0000_0213; // 0000_0000_0000_0000_0000_0100_0001_0011
        // ram[10] = 32'h0000_0013; // 0000_0000_0000_0000_0000_0000_0001_0011
        // ram[11] = 32'h0000_0013; // 0000_0000_0000_0000_0000_0000_0001_0011
        // // LOOP_J
        // ram[12] = 32'h04a2_0a63; // 0000_0100_1010_0010_0000_0110_0110_0011
        // ram[13] = 32'h0000_0293; // 0000_0000_0000_0000_0000_0101_0001_0011
        // ram[14] = 32'h0000_0013; // 0000_0000_0000_0000_0000_0000_0001_0011
        // ram[15] = 32'h0000_0013; // 0000_0000_0000_0000_0000_0000_0001_0011
        // // LOOP_K
        // ram[16] = 32'h02a2_8a63; // 0000_0010_1010_0010_1000_1010_0110_0011
        // ram[17] = 32'h00a1_85b3; // 0000_0000_1010_0011_0000_0101_1011_0011
        // ram[18] = 32'h0055_85b3; // 0000_0000_0101_0101_1000_0101_1011_0011
        // ram[19] = 32'h0025_9593; // 0000_0000_1001_0101_1010_0101_1011_0011
        // ram[20] = 32'h0005_a603; // 0000_0000_0000_0101_1010_0110_0000_0011
        // ram[21] = 32'h00a2_85b3; // 0000_0000_1010_0010_1000_0101_1011_0011
        // ram[22] = 32'h0045_85b3; // 0000_0000_0100_0101_1010_0101_1011_0011
        // ram[23] = 32'h0025_9593; // 0000_0000_1001_0101_1010_0101_1011_0011
        // ram[24] = 32'h0005_a683; // 0000_0000_0000_0101_1010_0110_1000_0011
        // ram[25] = 32'h00d6_06b3; // 0000_0000_1101_0110_0000_0110_1011_0011
        // ram[26] = 32'h00e6_8733; // 0000_0000_1110_0110_1010_0111_0011_0011
        // ram[27] = 32'h0012_8293; // 0000_0000_0001_0010_1000_0101_0001_0011
        // ram[28] = 32'hfc00_08e3; // 1111_1100_0000_0000_0000_1000_1110_0011
        // // LOOP_K_DONE
        // ram[29] = 32'h0000_0013;
        // ram[30] = 32'h0000_0013;
        // ram[31] = 32'h0012_0213; // 0000_0000_0001_0010_0000_0101_0001_0011
        // ram[32] = 32'hfa00_08e3; // 1111_1010_0000_0000_0011_1100_1110_0011
        // // LOOP_J_DONE
        // ram[33] = 32'h0000_0013;
        // ram[34] = 32'h0000_0013;
        // ram[35] = 32'h0011_8193; // 0000_0000_0001_0001_1000_0011_0001_0011
        // ram[36] = 32'hf800_08e3; // 1111_1010_0000_0000_0000_0000_1110_0011
        // // LOOP_I_DONE
        // ram[37] = 32'h0000_8067; // 0000_0000_0000_0000_1000_0000_0110_0111
        // // DONE
        // ram[38] = 32'h0000_0013; // 0000_0000_0000_0000_0000_0000_0001_0011
        // ram[39] = 32'h0000_0013; // 0000_0000_0000_0000_0000_0000_0001_0011


    // end
    
    
    always @(posedge clk) begin
        if (write_enable) begin
            ram[word_address] <= write_data;
        end 
    end
    
    assign read_data = ram[word_address];
    // assign next_read_data = ram[word_address + 1];
    // assign pc_inc = byte_address + 4;
endmodule
