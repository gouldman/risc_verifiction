package tb_pkg;
    import uvm_pkg::*; 
    `include "uvm_macros.svh"
    `include "alu_transaction.sv"
    `include "alu_in_monitor.sv"
    `include "alu_driver.sv"
    `include "alu_env.sv"
endpackage