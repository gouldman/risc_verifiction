// You can insert code here by setting file_header_inc in file execute_common.tpl

//=============================================================================
// Project  : generated_execute_tb
//
// File Name: forward_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Wed Nov 12 19:32:24 2025
//=============================================================================
// Description: Package for agent forward
//=============================================================================

package forward_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;


  `include "forward_forward_tx.sv"
  `include "forward_config.sv"
  `include "forward_driver.sv"
  `include "forward_monitor.sv"
  `include "forward_sequencer.sv"
  `include "forward_coverage.sv"
  `include "forward_agent.sv"
  `include "forward_seq_lib.sv"

endpackage : forward_pkg
